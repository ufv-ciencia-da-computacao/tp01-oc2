module shiftLeft(	input [63:0] dataIn,
						input [63:0] dataOut);


						
endmodule
