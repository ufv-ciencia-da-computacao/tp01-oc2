module immGenerator(	input [31:0] instruction,
							output [63:0] immediate);

		

endmodule
