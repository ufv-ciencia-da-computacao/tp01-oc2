module aluControl();

endmodule
